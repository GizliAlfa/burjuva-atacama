module aio20(
	AIO20_SPI_CLK_IN,
	AIO20_SPI_CLK_OUT,
	AIO20_SPI_MOSI_IN,
	AIO20_SPI_MOSI_OUT,
	AIO20_SPI_MISO_IN,
	AIO20_SPI_MISO_OUT,
	AIO20_SPI_NSS_IN,
	AIO20_SPI_NSS_OUT,
	AIO20_SPI_INT_IN,
	AIO20_SPI_INT_OUT,
	AIO20_CNVT_IN,
	AIO20_CNVT_OUT
);

input AIO20_SPI_CLK_IN; 
output AIO20_SPI_CLK_OUT; 
input AIO20_SPI_MOSI_IN; 
output AIO20_SPI_MOSI_OUT; 
input AIO20_SPI_MISO_IN; 
output AIO20_SPI_MISO_OUT; 
input AIO20_SPI_NSS_IN; 
output AIO20_SPI_NSS_OUT; 
input AIO20_SPI_INT_IN; 
output AIO20_SPI_INT_OUT; 
input AIO20_CNVT_IN; 
output AIO20_CNVT_OUT; 



assign AIO20_SPI_CLK_OUT = AIO20_SPI_NSS_IN == 0 ? AIO20_SPI_CLK_IN : 0;
assign AIO20_SPI_MOSI_OUT = AIO20_SPI_NSS_IN == 0 ? AIO20_SPI_MOSI_IN : 0;
assign AIO20_SPI_MISO_OUT = AIO20_SPI_NSS_IN == 0 ? AIO20_SPI_MISO_IN : 0;
assign AIO20_SPI_NSS_OUT = AIO20_SPI_NSS_IN;
assign AIO20_SPI_INT_OUT = AIO20_SPI_INT_IN;
assign AIO20_CNVT_OUT = AIO20_CNVT_IN;


endmodule
