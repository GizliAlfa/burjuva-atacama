module io16(
	IO16_SPI_CLK_IN,
	IO16_SPI_CLK_OUT,
	IO16_SPI_MOSI_IN,
	IO16_SPI_MOSI_OUT,
	IO16_SPI_MISO_IN,
	IO16_SPI_MISO_OUT,
	IO16_SPI_NSS_IN,
	IO16_SPI_NSS_OUT,
	IO16_SPI_INT_IN,
	IO16_SPI_INT_OUT
);

input IO16_SPI_CLK_IN; 
output IO16_SPI_CLK_OUT; 
input IO16_SPI_MOSI_IN; 
output IO16_SPI_MOSI_OUT; 
input IO16_SPI_MISO_IN; 
output IO16_SPI_MISO_OUT; 
input IO16_SPI_NSS_IN; 
output IO16_SPI_NSS_OUT; 
input IO16_SPI_INT_IN; 
output IO16_SPI_INT_OUT; 



assign IO16_SPI_CLK_OUT = IO16_SPI_CLK_IN;
assign IO16_SPI_MOSI_OUT = IO16_SPI_MOSI_IN;
assign IO16_SPI_MISO_OUT = IO16_SPI_MISO_IN;
assign IO16_SPI_NSS_OUT = IO16_SPI_NSS_IN;
assign IO16_SPI_INT_OUT = IO16_SPI_INT_IN;


endmodule
