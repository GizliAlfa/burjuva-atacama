module fpga(
	FPGA_SPI_CLK_IN,
	FPGA_SPI_CLK_OUT,
	FPGA_SPI_MOSI_IN,
	FPGA_SPI_MOSI_OUT,
	FPGA_SPI_MISO_IN,
	FPGA_SPI_MISO_OUT,
	FPGA_SPI_NSS_IN,
	FPGA_SPI_NSS_OUT,
	FPGA_SPI_INT_IN,
	FPGA_SPI_INT_OUT,
	FPGA_CRESET_IN,
	FPGA_CRESET_OUT,
	FPGA_CDONE_IN,
	FPGA_CDONE_OUT
);

input FPGA_SPI_CLK_IN; 
output FPGA_SPI_CLK_OUT; 
input FPGA_SPI_MOSI_IN; 
output FPGA_SPI_MOSI_OUT; 
input FPGA_SPI_MISO_IN; 
output FPGA_SPI_MISO_OUT; 
input FPGA_SPI_NSS_IN; 
output FPGA_SPI_NSS_OUT; 
input FPGA_SPI_INT_IN; 
output FPGA_SPI_INT_OUT; 
input FPGA_CRESET_IN; 
output FPGA_CRESET_OUT; 
input FPGA_CDONE_IN; 
output FPGA_CDONE_OUT; 



assign FPGA_SPI_CLK_OUT = FPGA_SPI_NSS_IN == 0 ? FPGA_SPI_CLK_IN : 0;
assign FPGA_SPI_MOSI_OUT = FPGA_SPI_NSS_IN == 0 ? FPGA_SPI_MOSI_IN : 0;
assign FPGA_SPI_MISO_OUT = FPGA_SPI_NSS_IN == 0 ? FPGA_SPI_MISO_IN : 0;
assign FPGA_SPI_NSS_OUT = FPGA_SPI_NSS_IN;
assign FPGA_SPI_INT_OUT = FPGA_SPI_INT_IN;
assign FPGA_CRESET_OUT = FPGA_CRESET_IN;
assign FPGA_CDONE_OUT = FPGA_CDONE_IN;


endmodule
